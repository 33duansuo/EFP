`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SEU
// Engineer: Renjun Duan
// 
// Create Date: 2024/12/15 16:46:45
// Design Name: 
// Module Name: decimal_to_efp8
// Project Name: 
// Target Devices: decimal_to_efp8
// Tool Versions: vivado 2023.2
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module decimal_to_efp(
    input [31:0] decimal_input,    // 32λ����
    input clk,
    input rst,
    input button,
    output reg [7:0] efp_output    // ���8λEFP��ʾ
);

// ���ұ�16λʮ��������8λEFP��ӳ�䣩
reg [31:0] lut [0:127];  // ���ұ��С128����Ҫ�����ұ��ʵ�����ݣ�

// �����ź�
reg [31:0] receive;
reg [7:0] i;  // ѭ��������
reg flag_1=0;  // ������־λ

// ���ұ�ĳ�ʼ����ʾ����ʼ����ֻ����һ���֣�ʵ��Ӧ����ʵ�ʲ��ұ���д��
initial begin
    lut[0] = 32'h00000078;    // Example: 0 -> 8'b00000000
    lut[1] = 32'h00000085;    // Example: 1 -> 8'b00000001
    lut[2] = 32'h00000093;    // Example: 2 -> 8'b00000010
    lut[3] = 32'h00000101;    // Example: 3 -> 8'b00000011
    lut[4] = 32'h00000110;    // Example: 4 -> 8'b00000100
    lut[5] = 32'h00000120;    // Example: 5 -> 8'b00000101
    lut[6] = 32'h00000131;    // Example: 6 -> 8'b00000110
    lut[7] = 32'h00000143;    // Example: 7 -> 8'b00000111
    lut[8] = 32'h00000156;    // Example: 8 -> 8'b00001000
    lut[9] = 32'h00000170;    // Example: 9 -> 8'b00001001
    lut[10] = 32'h00000186;   // Example: 10 -> 8'b00001010
    lut[11] = 32'h00000203;   // Example: 11 -> 8'b00001011
    lut[12] = 32'h00000221;   // Example: 12 -> 8'b00001100
    lut[13] = 32'h00000241;   // Example: 13 -> 8'b00001101
    lut[14] = 32'h00000263;   // Example: 14 -> 8'b00001110
    lut[15] = 32'h00000287;   // Example: 15 -> 8'b00001111
    lut[16] = 32'h00000312;   // Example: 16 -> 8'b00010000
    lut[17] = 32'h00000341;   // Example: 17 -> 8'b00010001
    lut[18] = 32'h00000372;   // Example: 18 -> 8'b00010010
    lut[19] = 32'h00000405;   // Example: 19 -> 8'b00010011
    lut[20] = 32'h00000442;   // Example: 20 -> 8'b00010100
    lut[21] = 32'h00000482;   // Example: 21 -> 8'b00010101
    lut[22] = 32'h00000526;   // Example: 22 -> 8'b00010110
    lut[23] = 32'h00000573;   // Example: 23 -> 8'b00010111
    lut[24] = 32'h00000625;   // Example: 24 -> 8'b00011000
    lut[25] = 32'h00000682;   // Example: 25 -> 8'b00011001
    lut[26] = 32'h00000743;   // Example: 26 -> 8'b00011010
    lut[27] = 32'h00000811;   // Example: 27 -> 8'b00011011
    lut[28] = 32'h00000884;   // Example: 28 -> 8'b00011100
    lut[29] = 32'h00000964;   // Example: 29 -> 8'b00011101
    lut[30] = 32'h00001051;   // Example: 30 -> 8'b00011110
    lut[31] = 32'h00001146;   // Example: 31 -> 8'b00011111
    lut[32] = 32'h00001250;   // Example: 32 -> 8'b00100000
    lut[33] = 32'h00001363;   // Example: 33 -> 8'b00100001
    lut[34] = 32'h00001487;   // Example: 34 -> 8'b00100010
    lut[35] = 32'h00001621;   // Example: 35 -> 8'b00100011
    lut[36] = 32'h00001768;   // Example: 36 -> 8'b00100100
    lut[37] = 32'h00001928;   // Example: 37 -> 8'b00100101
    lut[38] = 32'h00002102;   // Example: 38 -> 8'b00100110
    lut[39] = 32'h00002293;   // Example: 39 -> 8'b00100111
    lut[40] = 32'h00002500;   // Example: 40 -> 8'b00101000
    lut[41] = 32'h00002726;   // Example: 41 -> 8'b00101001
    lut[42] = 32'h00002973;   // Example: 42 -> 8'b00101010
    lut[43] = 32'h00003242;   // Example: 43 -> 8'b00101011
    lut[44] = 32'h00003536;   // Example: 44 -> 8'b00101100
    lut[45] = 32'h00003856;   // Example: 45 -> 8'b00101101
    lut[46] = 32'h00004204;   // Example: 46 -> 8'b00101110
    lut[47] = 32'h00004585;   // Example: 47 -> 8'b00101111
    lut[48] = 32'h00005000;   // Example: 48 -> 8'b00110000
    lut[49] = 32'h00005453;   // Example: 49 -> 8'b00110001
    lut[50] = 32'h00005946;   // Example: 50 -> 8'b00110010
    lut[51] = 32'h00006484;   // Example: 51 -> 8'b00110011
    lut[52] = 32'h00007071;   // Example: 52 -> 8'b00110100
    lut[53] = 32'h00007711;   // Example: 53 -> 8'b00110101
    lut[54] = 32'h00008409;   // Example: 54 -> 8'b00110110
    lut[55] = 32'h00009170;   // Example: 55 -> 8'b00110111
    lut[56] = 32'h00010000;   // Example: 56 -> 8'b00111000
    lut[57] = 32'h00010905;   // Example: 57 -> 8'b00111001
    lut[58] = 32'h00011892;   // Example: 58 -> 8'b00111010
    lut[59] = 32'h00012968;   // Example: 59 -> 8'b00111011
    lut[60] = 32'h00014142;   // Example: 60 -> 8'b00111100
    lut[61] = 32'h00015422;   // Example: 61 -> 8'b00111101
    lut[62] = 32'h00016818;   // Example: 62 -> 8'b00111110
    lut[63] = 32'h00018340;   // Example: 63 -> 8'b00111111
    lut[64] = 32'h00020000;   // Example: 64 -> 8'b01000000
    lut[65] = 32'h00021810;   // Example: 65 -> 8'b01000001
    lut[66] = 32'h00023784;   // Example: 66 -> 8'b01000010
    lut[67] = 32'h00025937;   // Example: 67 -> 8'b01000011
    lut[68] = 32'h00028284;   // Example: 68 -> 8'b01000100
    lut[69] = 32'h00030844;   // Example: 69 -> 8'b01000101
    lut[70] = 32'h00033636;   // Example: 70 -> 8'b01000110
    lut[71] = 32'h00036680;   // Example: 71 -> 8'b01000111
    lut[72] = 32'h00040000;   // Example: 72 -> 8'b01001000
    lut[73] = 32'h00043620;   // Example: 73 -> 8'b01001001
    lut[74] = 32'h00047568;   // Example: 74 -> 8'b01001010
    lut[75] = 32'h00051874;   // Example: 75 -> 8'b01001011
    lut[76] = 32'h00056569;   // Example: 76 -> 8'b01001100
    lut[77] = 32'h00061688;   // Example: 77 -> 8'b01001101
    lut[78] = 32'h00067272;   // Example: 78 -> 8'b01001110
    lut[79] = 32'h00073360;   // Example: 79 -> 8'b01001111
    lut[80] = 32'h00080000;   // Example: 80 -> 8'b01010000    
    lut[81] = 32'h00087241;   // Example: 81 -> 8'b01010001
    lut[82] = 32'h00095137;   // Example: 82 -> 8'b01010010
    lut[83] = 32'h00103747;   // Example: 83 -> 8'b01010011
    lut[84] = 32'h00113137;   // Example: 84 -> 8'b01010100
    lut[85] = 32'h00123377;   // Example: 85 -> 8'b01010101
    lut[86] = 32'h00134543;   // Example: 86 -> 8'b01010110
    lut[87] = 32'h00146721;   // Example: 87 -> 8'b01010111
    lut[88] = 32'h00160000;   // Example: 88 -> 8'b01011000
    lut[89] = 32'h00174481;   // Example: 89 -> 8'b01011001
    lut[90] = 32'h00190273;   // Example: 90 -> 8'b01011010
    lut[91] = 32'h00207494;   // Example: 91 -> 8'b01011011
    lut[92] = 32'h00226274;   // Example: 92 -> 8'b01011100
    lut[93] = 32'h00246754;   // Example: 93 -> 8'b01011101
    lut[94] = 32'h00269087;   // Example: 94 -> 8'b01011110
    lut[95] = 32'h00293441;   // Example: 95 -> 8'b01011111
    lut[96] = 32'h00320000;   // Example: 96 -> 8'b01100000
    lut[97] = 32'h00348962;   // Example: 97 -> 8'b01100001
    lut[98] = 32'h00380546;   // Example: 98 -> 8'b01100010
    lut[99] = 32'h00414989;   // Example: 99 -> 8'b01100011
    lut[100] = 32'h00452548;  // Example: 100 -> 8'b01100100
    lut[101] = 32'h00493517;  // Example: 101 -> 8'b01100101
    lut[102] = 32'h00538174;  // Example: 102 -> 8'b01100110
    lut[103] = 32'h00586883;  // Example: 103 -> 8'b01100111
    lut[104] = 32'h00640000;  // Example: 104 -> 8'b01101000
    lut[105] = 32'h00697925;  // Example: 105 -> 8'b01101001
    lut[106] = 32'h00761093;  // Example: 106 -> 8'b01101010
    lut[107] = 32'h00829977;  // Example: 107 -> 8'b01101011
    lut[108] = 32'h00905097;  // Example: 108 -> 8'b01101100
    lut[109] = 32'h00987015;  // Example: 109 -> 8'b01101101
    lut[110] = 32'h01076347;  // Example: 110 -> 8'b01101110    
    lut[111] = 32'h01173765;  // Example: 111 -> 8'b01101111
    lut[112] = 32'h01280000;  // Example: 112 -> 8'b01110000
    lut[113] = 32'h01395850;  // Example: 113 -> 8'b01110001
    lut[114] = 32'h01522185;  // Example: 114 -> 8'b01110010
    lut[115] = 32'h01659955;  // Example: 115 -> 8'b01110011
    lut[116] = 32'h01810193;  // Example: 116 -> 8'b01110100
    lut[117] = 32'h01974030;  // Example: 117 -> 8'b01110101
    lut[118] = 32'h02152695;  // Example: 118 -> 8'b01110110
    lut[119] = 32'h02347530;  // Example: 119 -> 8'b01110111
    lut[120] = 32'h02560000;  // Example: 120 -> 8'b01111000
    lut[121] = 32'h02791700;  // Example: 121 -> 8'b01111001
    lut[122] = 32'h03044370;  // Example: 122 -> 8'b01111010
    lut[123] = 32'h03319909;  // Example: 123 -> 8'b01111011
    lut[124] = 32'h03620387;  // Example: 124 -> 8'b01111100
    lut[125] = 32'h03948060;  // Example: 125 -> 8'b01111101
    lut[126] = 32'h04305390;  // Example: 126 -> 8'b01111110
    lut[127] = 32'h04695061;  // Example: 127 -> 8'b01111111
    // Add other LUT entries as needed...
end

always @(posedge clk) begin
    receive<=decimal_input;
    if (rst) begin
        efp_output <= 8'h00;  // �������
        i <= 0;               // ��������
    end else if (button) begin
        // ��ʼ�����
        efp_output <= 8'h00;
        // �������(���⴦��)
         if (decimal_input[28] == 1'b1) begin
            flag_1 = 1;  // �������λΪ������־,������<=���������Ÿ�ֵ����Ӱ������ĸ�ֵ
            receive[31:28]=0;      // ȥ��������־λ
        end
        

        // �������ұ��ҵ����ʵ�����
        for (i = 0; i < 127; i = i + 1) begin
            if(receive==0)begin
                efp_output <= 8'h00;// 0�������ѭ��
                i = 127;// ǿ������ѭ��
            end
            else if (receive >= lut[i] && receive < lut[i+1]) begin
                efp_output <= i;  // ��������ֵ
                i = 127;          // ǿ������ѭ��
            end
        end
        if  (flag_1 == 1) begin
            efp_output[7]<= 1;  // �������
        end

    end
end


endmodule
