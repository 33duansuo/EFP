module efp8_to_decimal(
    input clk,            // ʱ���ź�
    input [2:0]E,
    input [2:0]M,
    input [7:0] efp8,       // ����� EFP8 ����
    output reg [51:0] decimal_value // �����ʮ���ƽ��������Ϊ 52 λ���
);
//     // �ڲ��źŶ���
//     reg sign;
//     reg [3:0] exponent_bits;
//     reg [2:0] mantissa_bits;
//     reg [3:0] exponent;
//     integer  mantissa;
//     reg [31:0] temp;
//     parameter BIAS1 = 4'd15;
//     parameter BIAS = 4'd7;


// always @(posedge clk) begin
//     if(E == 4 && M == 3) begin
//         // ��ȡ����λ��ָ��λ��β��λ
//         sign = efp8[7];
//         exponent_bits = efp8[6:3];
//         mantissa_bits = efp8[2:0];

//         // ��ʼ�����
//         decimal_value = 52'd0_00;
//         // ��������ֵ���
//         if (efp8 == 8'b00000000) begin
//             decimal_value = 52'd0_00; /_00/ ����ȫ��
//         end else if (efp8 == 8'b10000000) begin
//             decimal_value = 52'h0_0FFFF_00FFFF; // ��ʾ������
//         end else begin
//             // ����ָ����ȥ��ƫ��ֵ
//             exponent = exponent_bits - BIAS;

//             // ����β��ֵ
//             mantissa = mantissa_bits;

//             // ��������ֵ (-1)^sign * (2^exponent) * (2^(mantissa/8))
//             temp = 2.0 ** (mantissa/8.0); // ���� 2^(mantissa / 8) �ȼ������� 3 λ
//             if (sign == 1'b0) begin
//                 decimal_value = 100000*(temp*2**(exponent)); // ��ֵ
//             end else begin
//                 decimal_value = -100000*(temp*2**(exponent)); // ��ֵ
//             end
//         end
//     end
//     if(E == 5 && M == 2) begin
//         // ��ȡ����λ��ָ��λ��β��λ
//         sign = efp8[7];
//         exponent_bits = efp8[6:2];
//         mantissa_bits = efp8[1:0];

//         // ��ʼ�����
//         decimal_value = 52'd0_00;
//         // ��������ֵ���
//         if (efp8 == 8'b00000000) begin
//             decimal_value = 52'd0_00; /_00/ ����ȫ��
//         end else if (efp8 == 8'b10000000) begin
//             decimal_value = 52'h0_0FFFF_00FFFF; // ��ʾ������
//         end else begin
//             // ����ָ����ȥ��ƫ��ֵ
//             exponent = exponent_bits - BIAS1;

//             // ����β��ֵ
//             mantissa = mantissa_bits;

//             // ��������ֵ (-1)^sign * (2^exponent) * (2^(mantissa/8))
//             temp = (2 ** mantissa)/4; // ���� 2^(mantissa / 8) �ȼ������� 3 λ
//             if (sign == 1'b0) begin
//                 decimal_value = 100000*(temp*2**(exponent)); // ��ֵ
//             end else begin
//                 decimal_value = -100000*(temp*2**(exponent)); // ��ֵ
//             end
//         end
//     end
// end
reg [51:0] lutE5M2 [0:127];  
reg [51:0] lutE4M3 [0:127];  
initial begin
    lutE4M3[0] = 52'h0_000000_000078;    // Example: 0 -> 8'b00000000
    lutE4M3[1] = 52'h0_000000_000085;    // Example: 1 -> 8'b00000001
    lutE4M3[2] = 52'h0_000000_000093;    // Example: 2 -> 8'b00000010
    lutE4M3[3] = 52'h0_000000_000101;    // Example: 3 -> 8'b00000011
    lutE4M3[4] = 52'h0_000000_000110;    // Example: 4 -> 8'b00000100
    lutE4M3[5] = 52'h0_000000_000120;    // Example: 5 -> 8'b00000101
    lutE4M3[6] = 52'h0_000000_000131;    // Example: 6 -> 8'b00000110
    lutE4M3[7] = 52'h0_000000_000143;    // Example: 7 -> 8'b00000111
    lutE4M3[8] = 52'h0_000000_000156;    // Example: 8 -> 8'b00001000
    lutE4M3[9] = 52'h0_000000_000170;    // Example: 9 -> 8'b00001001
    lutE4M3[10] = 52'h0_000000_000186;   // Example: 10 -> 8'b00001010
    lutE4M3[11] = 52'h0_000000_000203;   // Example: 11 -> 8'b00001011
    lutE4M3[12] = 52'h0_000000_000221;   // Example: 12 -> 8'b00001100
    lutE4M3[13] = 52'h0_000000_000241;   // Example: 13 -> 8'b00001101
    lutE4M3[14] = 52'h0_000000_000263;   // Example: 14 -> 8'b00001110
    lutE4M3[15] = 52'h0_000000_000287;   // Example: 15 -> 8'b00001111
    lutE4M3[16] = 52'h0_000000_000312;   // Example: 16 -> 8'b00010000
    lutE4M3[17] = 52'h0_000000_000341;   // Example: 17 -> 8'b00010001
    lutE4M3[18] = 52'h0_000000_000372;   // Example: 18 -> 8'b00010010
    lutE4M3[19] = 52'h0_000000_000405;   // Example: 19 -> 8'b00010011
    lutE4M3[20] = 52'h0_000000_000442;   // Example: 20 -> 8'b00010100
    lutE4M3[21] = 52'h0_000000_000482;   // Example: 21 -> 8'b00010101
    lutE4M3[22] = 52'h0_000000_000526;   // Example: 22 -> 8'b00010110
    lutE4M3[23] = 52'h0_000000_000573;   // Example: 23 -> 8'b00010111
    lutE4M3[24] = 52'h0_000000_000625;   // Example: 24 -> 8'b00011000
    lutE4M3[25] = 52'h0_000000_000682;   // Example: 25 -> 8'b00011001
    lutE4M3[26] = 52'h0_000000_000743;   // Example: 26 -> 8'b00011010
    lutE4M3[27] = 52'h0_000000_000811;   // Example: 27 -> 8'b00011011
    lutE4M3[28] = 52'h0_000000_000884;   // Example: 28 -> 8'b00011100
    lutE4M3[29] = 52'h0_000000_000964;   // Example: 29 -> 8'b00011101
    lutE4M3[30] = 52'h0_000000_001051;   // Example: 30 -> 8'b00011110
    lutE4M3[31] = 52'h0_000000_001146;   // Example: 31 -> 8'b00011111
    lutE4M3[32] = 52'h0_000000_001250;   // Example: 32 -> 8'b00100000
    lutE4M3[33] = 52'h0_000000_001363;   // Example: 33 -> 8'b00100001
    lutE4M3[34] = 52'h0_000000_001487;   // Example: 34 -> 8'b00100010
    lutE4M3[35] = 52'h0_000000_001621;   // Example: 35 -> 8'b00100011
    lutE4M3[36] = 52'h0_000000_001768;   // Example: 36 -> 8'b00100100
    lutE4M3[37] = 52'h0_000000_001928;   // Example: 37 -> 8'b00100101
    lutE4M3[38] = 52'h0_000000_002102;   // Example: 38 -> 8'b00100110
    lutE4M3[39] = 52'h0_000000_002293;   // Example: 39 -> 8'b00100111
    lutE4M3[40] = 52'h0_000000_002500;   // Example: 40 -> 8'b00101000
    lutE4M3[41] = 52'h0_000000_002726;   // Example: 41 -> 8'b00101001
    lutE4M3[42] = 52'h0_000000_002973;   // Example: 42 -> 8'b00101010
    lutE4M3[43] = 52'h0_000000_003242;   // Example: 43 -> 8'b00101011
    lutE4M3[44] = 52'h0_000000_003536;   // Example: 44 -> 8'b00101100
    lutE4M3[45] = 52'h0_000000_003856;   // Example: 45 -> 8'b00101101
    lutE4M3[46] = 52'h0_000000_004204;   // Example: 46 -> 8'b00101110
    lutE4M3[47] = 52'h0_000000_004585;   // Example: 47 -> 8'b00101111
    lutE4M3[48] = 52'h0_000000_005000;   // Example: 48 -> 8'b00110000
    lutE4M3[49] = 52'h0_000000_005453;   // Example: 49 -> 8'b00110001
    lutE4M3[50] = 52'h0_000000_005946;   // Example: 50 -> 8'b00110010
    lutE4M3[51] = 52'h0_000000_006484;   // Example: 51 -> 8'b00110011
    lutE4M3[52] = 52'h0_000000_007071;   // Example: 52 -> 8'b00110100
    lutE4M3[53] = 52'h0_000000_007711;   // Example: 53 -> 8'b00110101
    lutE4M3[54] = 52'h0_000000_008409;   // Example: 54 -> 8'b00110110
    lutE4M3[55] = 52'h0_000000_009170;   // Example: 55 -> 8'b00110111
    lutE4M3[56] = 52'h0_000001_000000;   // Example: 56 -> 8'b00111000
    lutE4M3[57] = 52'h0_000001_000905;   // Example: 57 -> 8'b00111001
    lutE4M3[58] = 52'h0_000001_001892;   // Example: 58 -> 8'b00111010
    lutE4M3[59] = 52'h0_000001_002968;   // Example: 59 -> 8'b00111011
    lutE4M3[60] = 52'h0_000001_004142;   // Example: 60 -> 8'b00111100
    lutE4M3[61] = 52'h0_000001_005422;   // Example: 61 -> 8'b00111101
    lutE4M3[62] = 52'h0_000001_006818;   // Example: 62 -> 8'b00111110
    lutE4M3[63] = 52'h0_000001_008340;   // Example: 63 -> 8'b00111111
    lutE4M3[64] = 52'h0_000002_000000;   // Example: 64 -> 8'b01000000
    lutE4M3[65] = 52'h0_000002_001810;   // Example: 65 -> 8'b01000001
    lutE4M3[66] = 52'h0_000002_003784;   // Example: 66 -> 8'b01000010
    lutE4M3[67] = 52'h0_000002_005937;   // Example: 67 -> 8'b01000011
    lutE4M3[68] = 52'h0_000002_008284;   // Example: 68 -> 8'b01000100
    lutE4M3[69] = 52'h0_000003_000844;   // Example: 69 -> 8'b01000101
    lutE4M3[70] = 52'h0_000003_003636;   // Example: 70 -> 8'b01000110
    lutE4M3[71] = 52'h0_000003_006680;   // Example: 71 -> 8'b01000111
    lutE4M3[72] = 52'h0_000004_000000;   // Example: 72 -> 8'b01001000
    lutE4M3[73] = 52'h0_000004_003620;   // Example: 73 -> 8'b01001001
    lutE4M3[74] = 52'h0_000004_007568;   // Example: 74 -> 8'b01001010
    lutE4M3[75] = 52'h0_000005_001874;   // Example: 75 -> 8'b01001011
    lutE4M3[76] = 52'h0_000005_006569;   // Example: 76 -> 8'b01001100
    lutE4M3[77] = 52'h0_000006_001688;   // Example: 77 -> 8'b01001101
    lutE4M3[78] = 52'h0_000006_007272;   // Example: 78 -> 8'b01001110
    lutE4M3[79] = 52'h0_000007_003360;   // Example: 79 -> 8'b01001111
    lutE4M3[80] = 52'h0_000008_000000;   // Example: 80 -> 8'b01010000    
    lutE4M3[81] = 52'h0_000008_007241;   // Example: 81 -> 8'b01010001
    lutE4M3[82] = 52'h0_000009_005137;   // Example: 82 -> 8'b01010010
    lutE4M3[83] = 52'h0_000010_003747;   // Example: 83 -> 8'b01010011
    lutE4M3[84] = 52'h0_000011_003137;   // Example: 84 -> 8'b01010100
    lutE4M3[85] = 52'h0_000012_003377;   // Example: 85 -> 8'b01010101
    lutE4M3[86] = 52'h0_000013_004543;   // Example: 86 -> 8'b01010110
    lutE4M3[87] = 52'h0_000014_006721;   // Example: 87 -> 8'b01010111
    lutE4M3[88] = 52'h0_000016_000000;   // Example: 88 -> 8'b01011000
    lutE4M3[89] = 52'h0_000017_004481;   // Example: 89 -> 8'b01011001
    lutE4M3[90] = 52'h0_000019_000273;   // Example: 90 -> 8'b01011010
    lutE4M3[91] = 52'h0_000020_007494;   // Example: 91 -> 8'b01011011
    lutE4M3[92] = 52'h0_000022_006274;   // Example: 92 -> 8'b01011100
    lutE4M3[93] = 52'h0_000024_006754;   // Example: 93 -> 8'b01011101
    lutE4M3[94] = 52'h0_000026_009087;   // Example: 94 -> 8'b01011110
    lutE4M3[95] = 52'h0_000029_003441;   // Example: 95 -> 8'b01011111
    lutE4M3[96] = 52'h0_000032_000000;   // Example: 96 -> 8'b01100000
    lutE4M3[97] = 52'h0_000034_008962;   // Example: 97 -> 8'b01100001
    lutE4M3[98] = 52'h0_000038_000546;   // Example: 98 -> 8'b01100010
    lutE4M3[99] = 52'h0_000041_004989;   // Example: 99 -> 8'b01100011
    lutE4M3[100] = 52'h0_000045_002548;  // Example: 100 -> 8'b01100100
    lutE4M3[101] = 52'h0_000049_003517;  // Example: 101 -> 8'b01100101
    lutE4M3[102] = 52'h0_000053_008174;  // Example: 102 -> 8'b01100110
    lutE4M3[103] = 52'h0_000058_006883;  // Example: 103 -> 8'b01100111
    lutE4M3[104] = 52'h0_000064_000000;  // Example: 104 -> 8'b01101000
    lutE4M3[105] = 52'h0_000069_007925;  // Example: 105 -> 8'b01101001
    lutE4M3[106] = 52'h0_000076_001093;  // Example: 106 -> 8'b01101010
    lutE4M3[107] = 52'h0_000082_009977;  // Example: 107 -> 8'b01101011
    lutE4M3[108] = 52'h0_000090_005097;  // Example: 108 -> 8'b01101100
    lutE4M3[109] = 52'h0_000098_007015;  // Example: 109 -> 8'b01101101
    lutE4M3[110] = 52'h0_000107_006347;  // Example: 110 -> 8'b01101110    
    lutE4M3[111] = 52'h0_000117_003765;  // Example: 111 -> 8'b01101111
    lutE4M3[112] = 52'h0_000128_000000;  // Example: 112 -> 8'b01110000
    lutE4M3[113] = 52'h0_000139_005850;  // Example: 113 -> 8'b01110001
    lutE4M3[114] = 52'h0_000152_002185;  // Example: 114 -> 8'b01110010
    lutE4M3[115] = 52'h0_000165_009955;  // Example: 115 -> 8'b01110011
    lutE4M3[116] = 52'h0_000181_000193;  // Example: 116 -> 8'b01110100
    lutE4M3[117] = 52'h0_000197_004030;  // Example: 117 -> 8'b01110101
    lutE4M3[118] = 52'h0_000215_002695;  // Example: 118 -> 8'b01110110
    lutE4M3[119] = 52'h0_000234_007530;  // Example: 119 -> 8'b01110111
    lutE4M3[120] = 52'h0_000256_000000;  // Example: 120 -> 8'b01111000
    lutE4M3[121] = 52'h0_000279_001700;  // Example: 121 -> 8'b01111001
    lutE4M3[122] = 52'h0_000304_004370;  // Example: 122 -> 8'b01111010
    lutE4M3[123] = 52'h0_000331_009909;  // Example: 123 -> 8'b01111011
    lutE4M3[124] = 52'h0_000362_000387;  // Example: 124 -> 8'b01111100
    lutE4M3[125] = 52'h0_000394_008060;  // Example: 125 -> 8'b01111101
    lutE4M3[126] = 52'h0_000430_005390;  // Example: 126 -> 8'b01111110
    lutE4M3[127] = 52'h0_000469_005061;  // Example: 127 -> 8'b01111111
    //E5M2
    lutE5M2[0]=52'h0_000000_000031;
    lutE5M2[1]=52'h0_000000_000036;
    lutE5M2[2]=52'h0_000000_000043;
    lutE5M2[3]=52'h0_000000_000051;
    lutE5M2[4]=52'h0_000000_000061;
    lutE5M2[5]=52'h0_000000_000073;
    lutE5M2[6]=52'h0_000000_000087;
    lutE5M2[7]=52'h0_000000_000103;
    lutE5M2[8]=52'h0_000000_000122;
    lutE5M2[9]=52'h0_000000_000145;
    lutE5M2[10]=52'h0_000000_000173;
    lutE5M2[11]=52'h0_000000_000205;
    lutE5M2[12]=52'h0_000000_000244;
    lutE5M2[13]=52'h0_000000_000290;
    lutE5M2[14]=52'h0_000000_000345;
    lutE5M2[15]=52'h0_000000_000411;
    lutE5M2[16]=52'h0_000000_000488;
    lutE5M2[17]=52'h0_000000_000581;
    lutE5M2[18]=52'h0_000000_000691;
    lutE5M2[19]=52'h0_000000_000821;
    lutE5M2[20]=52'h0_000000_000977;
    lutE5M2[21]=52'h0_000000_001161;
    lutE5M2[22]=52'h0_000000_001381;
    lutE5M2[23]=52'h0_000000_001642;
    lutE5M2[24]=52'h0_000000_001953;
    lutE5M2[25]=52'h0_000000_002323;
    lutE5M2[26]=52'h0_000000_002762;
    lutE5M2[27]=52'h0_000000_003285;
    lutE5M2[28]=52'h0_000000_003906;
    lutE5M2[29]=52'h0_000000_004645;
    lutE5M2[30]=52'h0_000000_005524;
    lutE5M2[31]=52'h0_000000_006570;
    lutE5M2[32]=52'h0_000000_007813;
    lutE5M2[33]=52'h0_000000_009291;
    lutE5M2[34]=52'h0_000000_011049;
    lutE5M2[35]=52'h0_000000_013139;
    lutE5M2[36]=52'h0_000000_015625;
    lutE5M2[37]=52'h0_000000_018581;
    lutE5M2[38]=52'h0_000000_022097;
    lutE5M2[39]=52'h0_000000_026278;
    lutE5M2[40]=52'h0_000000_031250;
    lutE5M2[41]=52'h0_000000_037163;
    lutE5M2[42]=52'h0_000000_044194;
    lutE5M2[43]=52'h0_000000_052556;
    lutE5M2[44]=52'h0_000000_062500;
    lutE5M2[45]=52'h0_000000_074325;
    lutE5M2[46]=52'h0_000000_088384;
    lutE5M2[47]=52'h0_000000_105112;
    lutE5M2[48]=52'h0_000000_125000;
    lutE5M2[49]=52'h0_000000_148651;
    lutE5M2[50]=52'h0_000000_176777;
    lutE5M2[51]=52'h0_000000_210224;
    lutE5M2[52]=52'h0_000000_250000;
    lutE5M2[53]=52'h0_000000_297302;
    lutE5M2[54]=52'h0_000000_353553;
    lutE5M2[55]=52'h0_000000_420448;
    lutE5M2[56]=52'h0_000000_500000;
    lutE5M2[57]=52'h0_000000_594603;
    lutE5M2[58]=52'h0_000000_707107;
    lutE5M2[59]=52'h0_000000_840896;
    lutE5M2[60]=52'h0_000001_000000;
    lutE5M2[61]=52'h0_000001_189207;
    lutE5M2[62]=52'h0_000001_414214;
    lutE5M2[63]=52'h0_000001_681793;
    lutE5M2[64]=52'h0_000002_000000;
    lutE5M2[65]=52'h0_000002_378414;
    lutE5M2[66]=52'h0_000002_828427;
    lutE5M2[67]=52'h0_000003_363586;
    lutE5M2[68]=52'h0_000004_000000;
    lutE5M2[69]=52'h0_000004_756828;
    lutE5M2[70]=52'h0_000005_656854;
    lutE5M2[71]=52'h0_000006_727171;
    lutE5M2[72]=52'h0_000008_000000;
    lutE5M2[73]=52'h0_000009_513657;
    lutE5M2[74]=52'h0_000011_313709;
    lutE5M2[75]=52'h0_000013_454343;
    lutE5M2[76]=52'h0_000016_000000;
    lutE5M2[77]=52'h0_000019_027313;
    lutE5M2[78]=52'h0_000022_627417;
    lutE5M2[79]=52'h0_000026_908685;
    lutE5M2[80]=52'h0_000032_000000;
    lutE5M2[81]=52'h0_000038_054628;
    lutE5M2[82]=52'h0_000045_254834;
    lutE5M2[83]=52'h0_000053_817371;
    lutE5M2[84]=52'h0_000064_000000;
    lutE5M2[85]=52'h0_000076_109255;
    lutE5M2[86]=52'h0_000090_509668;
    lutE5M2[87]=52'h0_000107_634741;
    lutE5M2[88]=52'h0_000128_000000;
    lutE5M2[89]=52'h0_000152_218511;
    lutE5M2[90]=52'h0_000181_019336;
    lutE5M2[91]=52'h0_000215_269482;
    lutE5M2[92]=52'h0_000256_000000;
    lutE5M2[93]=52'h0_000304_437021;
    lutE5M2[94]=52'h0_000362_038672;
    lutE5M2[95]=52'h0_000430_538965;
    lutE5M2[96]=52'h0_000512_000000;
    lutE5M2[97]=52'h0_000608_874043;
    lutE5M2[98]=52'h0_000724_077344;
    lutE5M2[99]=52'h0_000861_077929;
    lutE5M2[100]=52'h0_001024_000000;
    lutE5M2[101]=52'h0_001217_748094;
    lutE5M2[102]=52'h0_001448_154693;
    lutE5M2[103]=52'h0_001722_155861;
    lutE5M2[104]=52'h0_002048_000000;
    lutE5M2[105]=52'h0_002435_496173;
    lutE5M2[106]=52'h0_002896_309384;
    lutE5M2[107]=52'h0_003444_311717;
    lutE5M2[108]=52'h0_004096_000000;
    lutE5M2[109]=52'h0_004870_992347;
    lutE5M2[110]=52'h0_005792_618751;
    lutE5M2[111]=52'h0_006888_623429;
    lutE5M2[112]=52'h0_008192_000000;
    lutE5M2[113]=52'h0_009741_984692;
    lutE5M2[114]=52'h0_011585_237502;
    lutE5M2[115]=52'h0_013777_246892;
    lutE5M2[116]=52'h0_016384_000000;
    lutE5M2[117]=52'h0_019483_969423;
    lutE5M2[118]=52'h0_023170_475007;
    lutE5M2[119]=52'h0_027554_493708;
    lutE5M2[120]=52'h0_032768_000000;
    lutE5M2[121]=52'h0_038967_938673;
    lutE5M2[122]=52'h0_046340_950002;
    lutE5M2[123]=52'h0_055108_987506;
    lutE5M2[124]=52'h0_065536_000000;
    lutE5M2[125]=52'h0_077935_877508;
    lutE5M2[126]=52'h0_092681_900003;
    lutE5M2[127]=52'h0_110217_975118;

end

    always @ (posedge clk) begin
        if(E==4&&M==3) begin
        decimal_value <= lutE4M3[efp8];
        end 
        else if(E==5&&M==2) begin
        decimal_value <= lutE5M2[efp8];
        end 
    end

endmodule
